//---------------------------------------------------------
// ROM Module
//---------------------------------------------------------
module rom (
  input	 	[7:0]		data_in,
  output 	[7:0]		data_out
  );

endmodule
