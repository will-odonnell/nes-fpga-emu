//---------------------------------------------------------
// Input/Output Module
//---------------------------------------------------------
module io (
  input  	[7:0]		ctrl,
  input 	[15:0]		addr,
  inout  	[7:0]		data
  );

endmodule
