//---------------------------------------------------------
// MMC Module
//---------------------------------------------------------
module mmc (
  input  	[7:0]		ctrl,
  input 	[15:0]		addr,
  output	[7:0]		data
  );

endmodule
