//---------------------------------------------------------
// CPU module
//---------------------------------------------------------
module cpu(
  output 	[7:0]		ctrl,
  output 	[15:0]		addr,
  inout	 	[7:0]		data
  );

endmodule
